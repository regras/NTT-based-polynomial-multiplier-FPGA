library verilog;
use verilog.vl_types.all;
entity NTT_PolyMul_test is
end NTT_PolyMul_test;
